uno1_inst : uno1 PORT MAP (
		result	 => result_sig
	);
