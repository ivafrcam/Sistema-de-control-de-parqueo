dos4_inst : dos4 PORT MAP (
		result	 => result_sig
	);
