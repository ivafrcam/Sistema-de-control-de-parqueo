cuatro4_inst : cuatro4 PORT MAP (
		result	 => result_sig
	);
